----------------------------------------------------------------------
-- Digital Design 101 Lab Assignment 1 (Structural) - S22
-- LFDetector Structural Model
----------------------------------------------------------------------
-- Student First Name : Your First Name
-- Student Last Name : Your Last Name
-- Student ID : Your Student ID
----------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY NAND2 IS
   PORT (x: IN std_logic;
         y: IN std_logic;
         F: OUT std_logic);
END NAND2;  

ARCHITECTURE behav OF NAND2 IS
BEGIN
   PROCESS(x, y)
   BEGIN
      F <= NOT (x AND y) AFTER 1.4 ns; 
   END PROCESS;
END behav;
----------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY LFDetector_structural IS
   PORT (Fuel3, Fuel2, Fuel1, Fuel0: IN std_logic;
         FuelWarningLight: OUT std_logic);
END LFDetector_structural;

ARCHITECTURE Structural OF LFDetector_structural IS

-- DO NOT modify any signals, ports, or entities above this line
-- add your code below this line
-- you should be declaring and connecting components in this code
-- you should not use a PROCESS for lab 1s
-- use the appropriate library component(s) specified in the lab handout
-- add the appropriate internal signals & wire your design below
BEGIN
  FuelWarningLight <= NAND(NAND(NAND(Fuel3, Fuel3), NAND(Fuel2, Fuel2)), NAND(NAND(Fuel3, Fuel3), NAND(Fuel2, Fuel2)));
END Structural;